
module rom32(address, data_out);
  input  [31:0] address;
  output [31:0] data_out;
  reg    [31:0] data_out;

  parameter BASE_ADDRESS = 25'd0; // address that applies to this memory

  wire [6:0] mem_offset;
  wire address_select;

  assign mem_offset = address[7:2];  // drop 2 LSBs to get word offset

  assign address_select = (address[31:8] == BASE_ADDRESS);  // address decoding

  always @(address_select or mem_offset)

  begin
    if ((address % 4) != 0) $display($time, " rom32 error: unaligned address %d", address);
    if (address_select == 1)
    begin
      case (mem_offset)		
6'd0  : data_out = {32'b00011000000010100000000000000000};            //movi r5, #0 
6'd1  : data_out = {32'b00011000000011000001010111111000};            //movi r6, #5624
6'd2  : data_out = {32'b00011000000000100000000000000000};            //movi r1, #0
6'd3  : data_out = {32'b00011000000001000001010111111001};            //movi r2, #5625 
6'd4  : data_out = {32'b00011000000011100000000000000000};            //movi r7, #0 
6'd5  : data_out = {32'b00011000000100000000000000000000};            //movi r8, #0
6'd6  : data_out = {32'b00100000001010000000000010010110};            //mov.v v4, #150
6'd8  : data_out = {32'b01100001010011000000000000010101};            //beq r5, r6, desencriptar
6'd9  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd10  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd11  : data_out = {32'b01110000011100100000000000000000};            //load.v v9, r1
6'd12  : data_out = {32'b00000000000000000000000000000000};            //nop 
6'd13  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd14  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd15  : data_out = {32'b00010110011010010101000000000000};            //add.v v5, v9, v4
6'd16  : data_out = {32'b00000000000000000000000000000000};            //nop 
6'd17  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd18  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd19  : data_out = {32'b10000000101010100000000000000000};            //store.v v5, r2
6'd20  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd21  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd22  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd23  : data_out = {32'b10011000010000100000000000000001};            //addi r1, r1, #1
6'd24  : data_out = {32'b10011000100001000000000000000001};            //addi r2, r2, #1
6'd25  : data_out = {32'b10011001010010100000000000000001};            //addi r5, r5, #1
6'd26  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd27  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd28  : data_out = {32'b01100001110100011111111111101011};            //beq r7, r8, loop 
6'd29  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd31  : data_out = {32'b00011000000101000000000000000000};            //movi r10, #0 
6'd32  : data_out = {32'b00011000000101100001010111111000};            //movi r11, #5624
6'd33  : data_out = {32'b00011000000110000001010111111001};            //movi r12, #5625
6'd34  : data_out = {32'b00011000000110100010101111110010};            //movi r13, #11250
6'd36  : data_out = {32'b01100010100101100000000000010101};            //beq r10, r11, done
6'd37  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd38  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd39  : data_out = {32'b01110011001101000000000000000000};            //load.v v10, r12
6'd40  : data_out = {32'b00000000000000000000000000000000};            //nop 
6'd41  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd42  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd43  : data_out = {32'b10001110101010011011000000000000};            //sub.v v11, v10, v4
6'd44  : data_out = {32'b00000000000000000000000000000000};            //nop 
6'd45  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd46  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd47  : data_out = {32'b10000011011101100000000000000000};            //store.v v11, r13
6'd48  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd49  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd50  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd51  : data_out = {32'b10011011000110000000000000000001};            //addi r12, r12, #1
6'd52  : data_out = {32'b10011011010110100000000000000001};            //addi r13, r13, #1
6'd53  : data_out = {32'b10011010100101000000000000000001};            //addi r10, r10, #1
6'd54  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd55  : data_out = {32'b00000000000000000000000000000000};            //nop
6'd56  : data_out = {32'b01100001110100011111111111101011};            //beq r7, r8, loopDesencriptar 
6'd57  : data_out = {32'b00000000000000000000000000000000};            //nop
          default data_out = 32'h0000;
      endcase

   //   $display($time, " reading data: rom32[%h] => %h", address, data_out);

    end
  end
endmodule



