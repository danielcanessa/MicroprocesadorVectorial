//*** Instruction Set Definition in file "instruction_set.v" ***//
//*** TOP LEVEL MODULE ***//
module vemicry_module ( clock, reset, typ, data_read, data_write,
data_add, data_in_mem, memdataout, ID_VDF_VS_ADD, ID_VDF_VT_ADD, ID_VDF_VD_ADD,
ID_VDF_SHAMT, ID_VDF_OP, ID_VDF_FUNC, ID_VDF_IMM16, ID_VDF_INDEX, ID_EX_RS_VAL,
ID_EX_RT_VAL, pipe_stall, sbi_sig, sbi_add, sbi_val);

endmodule // Top Level VeMICry